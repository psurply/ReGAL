module top (
    input A,
    input B,
    output C,
    output D
);

assign C =
  (~A)
;

assign D =
  (~B)
;

endmodule
