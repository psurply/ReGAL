module top (
    input A,
    input B,
    output C
);

assign C =
  1
;

endmodule
